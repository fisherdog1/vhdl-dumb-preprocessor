�� 
 l i b r a r y   w o r k ;  
 	 u s e   w o r k . a d d r e s s _ m a t h . a l l ;  
  
 e n t i t y   u n i t _ t e s t s   i s  
 e n d   e n t i t y ;  
  
 a r c h i t e c t u r e   s i m   o f   u n i t _ t e s t s   i s  
 b e g i n  
 	 p r o c e s s  
 	 b e g i n  
 	 	 l o o p  
 	 	 	 r e p o r t   " m y _ f u n c t i o n ( 1 )   = =   2 "   s e v e r i t y   n o t e ;  
 	 	 	  
 	 	 	 i f   n o t   ( m y _ f u n c t i o n ( 1 )   = =   2 )   t h e n    
 	 	 	 	 r e p o r t   " F A I L "   s e v e r i t y   e r r o r ;  
 	 	 	 	 e x i t ;    
 	 	 	 e n d   i f ;  
 	 	 	  
 	 	 	 r e p o r t   " m y _ f u n c t i o n ( 3 )   = =   4 "   s e v e r i t y   n o t e ;  
 	 	 	  
 	 	 	 i f   n o t   ( m y _ f u n c t i o n ( 3 )   = =   4 )   t h e n    
 	 	 	 	 r e p o r t   " F A I L "   s e v e r i t y   e r r o r ;  
 	 	 	 	 e x i t ;    
 	 	 	 e n d   i f ;  
 	 	 	  
 	 	 	 a s s e r t   f a l s e   r e p o r t   " T e s t s   ! P A S S ! "   s e v e r i t y   f a i l u r e ;  
 	 	 e n d   l o o p ;  
  
 	 	 a s s e r t   f a l s e   r e p o r t   " T e s t s   ! F A I L ! "   s e v e r i t y   f a i l u r e ;  
 	 e n d   p r o c e s s ;  
 e n d   a r c h i t e c t u r e   s i m ;  
  
 