--snippets conditions
my_function(1) == 2
my_function(3) == 4
--endsnippets